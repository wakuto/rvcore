`ifndef RISCV_INSTR_H
`define RISCV_INSTR_H

`include "inst.sverilog"

`endif
